--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   11:32:42 08/21/2018
-- Design Name:   
-- Module Name:   C:/ProySisDigAva/HW2/HW2_tb.vhd
-- Project Name:  HW2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: HW2
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY HW2_tb IS
END HW2_tb;
 
ARCHITECTURE behavior OF HW2_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT HW2
    PORT(
         A : IN  std_logic;
         B : IN  std_logic;
         C : IN  std_logic;
         Y : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic := '0';
   signal B : std_logic := '0';
   signal C : std_logic := '0';

 	--Outputs
   signal Y : std_logic;
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: HW2 PORT MAP (
          A => A,
          B => B,
          C => C,
          Y => Y
        );

   -- Clock process definitions
--   <clock>_process :process
--   begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      --wait for <clock>_period*10;

      -- insert stimulus here 
		A <= '0'; B <= '0'; C <= '0'; wait for 100ns;
		A <= '0'; B <= '0'; C <= '1'; wait for 100ns;
		A <= '0'; B <= '1'; C <= '0'; wait for 100ns;
		A <= '0'; B <= '1'; C <= '1'; wait for 100ns;
		A <= '1'; B <= '0'; C <= '0'; wait for 100ns;
		A <= '1'; B <= '0'; C <= '1'; wait for 100ns;
		A <= '1'; B <= '1'; C <= '0'; wait for 100ns;
		A <= '1'; B <= '1'; C <= '1'; wait for 100ns;
      wait;
   end process;

END;
